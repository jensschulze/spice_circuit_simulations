psu simmons sds 800
.include ./lib/regulators.lib
v1 0 1 0 sin(0 12 50 0 0)
v2 2 0 0 sin(0 12 50 0 0)
rlast1 5 0 10k
rlast2 0 6 10k
d2 1 3 mod1
d3 2 3 mod1
d4 4 2 mod1
d5 4 1 mod1
c1 0 4 2200UF
c2 0 6 10UF
c3 0 6 0.1UF
c4 3 0 2200UF
c5 5 0 10UF
c6 5 0 0.1UF
X2 3 0 5 lm7805
X1 4 0 6 lm7905
d1 7 3 mod1
c7 7 0 220UF
.model mod1 d
.tran .5m 25m .1m
.save tran v(5) v(6)
.end
